../synth/binary.vhdl